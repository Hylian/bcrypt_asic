module sram ();


endmodule: sram
