module testbench;

   logic clk;

   bcrypt core(clk, , , );

endmodule: testbench
